module inst_memory_wrapper(



);



endmodule