module proc(



);








endmodule