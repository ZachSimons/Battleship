module memory_tester()



endmodule