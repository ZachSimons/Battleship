// Have two IPs (one for D-Memory and one for I-Memory)