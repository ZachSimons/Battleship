module eth_top (
    input  logic clk,
    input  logic rst_n,
    input  logic [31:0] data_in,
    input  logic        dval_in,
    output logic [31:0] data_out,
    output logic        dval_out
);


endmodule