module fetch(
    input branch
    input rti
    input interrupt


    input []


//Add one if making imem byte addressable


);



endmodule